**.subckt ampb vdd vss ip im o ib
*.iopin vdd
*.iopin vss
*.iopin ip
*.iopin im
*.iopin o
*.iopin ib
x1a ib ib vdd vdd p1_4
x2a x ib vdd vdd p1_4
x3a x ib vdd vdd p1_4
x3c __UNCONNECTED_PIN__0 net1 __UNCONNECTED_PIN__1 __UNCONNECTED_PIN__2 n1_4
x2c y __UNCONNECTED_PIN__3 vss vss n1_4
x2b __UNCONNECTED_PIN__4 ip x vdd p1_4
x3b __UNCONNECTED_PIN__5 im x vdd p1_4
x1 net5 net5 __UNCONNECTED_PIN__6 __UNCONNECTED_PIN__7 p1_4
x2 net5 __UNCONNECTED_PIN__8 net3 net3 n1_4
x3 net6 net5 __UNCONNECTED_PIN__9 __UNCONNECTED_PIN__10 p1_4
x4 net6 __UNCONNECTED_PIN__11 net4 net4 n1_4
**.ends

* expanding   symbol:  p1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_4.sch
.subckt p1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_2
xd D G X B p1_2
.ends


* expanding   symbol:  n1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_4.sch
.subckt n1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_2
xs X G S B n1_2
.ends


* expanding   symbol:  p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
