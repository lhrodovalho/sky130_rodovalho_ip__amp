**.subckt ampc_tb
iib_df ib_df GND {xib} 
cl_df o_df GND 'xc' m=1 
Xdut_df x_df cm o_df ib_df vdd_df GND ampc
vcm cm GND DC {xcm} 
ci_df in x_df 1T m=1
lf_df o_df x_df 1T m=1
vvdd_df vdd_df GND {xvdd} 
vin in cm DC 0 AC 1
iib_cm ib_cm GND {xib} 
cl_cm o_cm GND 'xc' m=1 
Xdut_cm x_cm in o_cm ib_cm vdd_cm GND ampc
ci_cm in x_cm 1T m=1
lf_cm o_cm x_cm 1T m=1
vvdd_cm vdd_cm GND {xvdd} 
iib_ps ib_ps GND {xib} 
cl_ps o_ps GND 'xc' m=1 
Xdut_ps x_ps cm o_ps ib_ps vdd_ps GND ampc
ci_ps cm x_ps 1T m=1
lf_ps o_ps x_ps 1T m=1
vvdd_ps vdd_ps GND DC {xvdd} AC 1 
**** begin user architecture code


* Include SkyWater sky130 device models
.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.param mc_mm_switch=0





.option gmin=1E-15
.control

  ac dec 10 1 1G
  let av_df = db(o_df)
  let ph_df = cphase(o_df)*180/(atan(1)*4)
  let av_cm = db(o_cm)
  let cmrr  = av_df-av_cm
  let av_ps = db(o_ps)
  let psrr  = av_df-av_ps

  plot av_df
  plot ph_df
  plot cmrr
  plot psrr

  meas ac av_1hz find av_df at=1
  meas ac cmrr_1hz find cmrr at=1
  meas ac psrr_1hz find cmrr at=1
  meas ac gbw when av_df=0
  meas ac pm find ph_df at=gbw

.endc




.param xvdd = 1.8
.param xcm  = 0.9
.param xib  = 100n
.param xc   = 1p


**** end user architecture code
**.ends

* expanding   symbol:  ampc.sym # of pins=6
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/ampc.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/ampc.sch
.subckt ampc  im  ip  o  ib  vdd  vss
*.iopin vdd
*.iopin vss
*.iopin ip
*.iopin im
*.iopin o
*.iopin ib
x1a ib ib vdd vdd p1_4
x2a x ib vdd vdd p1_4
x3a x ib vdd vdd p1_4
x3c z y vss vss n1_4
x2c y y vss vss n1_4
x2b y im x vdd p1_4
x3b z ip x vdd p1_4
x4a o ib vdd vdd p4_1
x4c o z vss vss n4_1
XC1 z o sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
.ends


* expanding   symbol:  p1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_4.sch
.subckt p1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_2
xd D G X B p1_2
.ends


* expanding   symbol:  n1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_4.sch
.subckt n1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_2
xs X G S B n1_2
.ends


* expanding   symbol:  p4_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p4_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p4_1.sch
.subckt p4_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p2_1
xr D G S B p2_1
.ends


* expanding   symbol:  n4_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n4_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n4_1.sch
.subckt n4_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n2_1
xl D G S B n2_1
.ends


* expanding   symbol:  p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  p2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p2_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p2_1.sch
.subckt p2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p1_1
xr D G S B p1_1
.ends


* expanding   symbol:  n2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n2_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n2_1.sch
.subckt n2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n1_1
xl D G S B n1_1
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/amp_tb/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
