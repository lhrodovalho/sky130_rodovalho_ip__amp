**.subckt ampc vdd vss ip im o ib
*.iopin vdd
*.iopin vss
*.iopin ip
*.iopin im
*.iopin o
*.iopin ib
x1a ib ib vdd vdd p1_4
x2a x ib vdd vdd p1_4
x3a x ib vdd vdd p1_4
x3c z y vss vss n1_4
x2c y y vss vss n1_4
x2b y im x vdd p1_4
x3b z ip x vdd p1_4
x4a o ib vdd vdd p4_1
x4c o z vss vss n4_1
XC1 z o sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
**.ends

* expanding   symbol:  p1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_4.sch
.subckt p1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_2
xd D G X B p1_2
.ends


* expanding   symbol:  n1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_4.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_4.sch
.subckt n1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_2
xs X G S B n1_2
.ends


* expanding   symbol:  p4_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p4_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p4_1.sch
.subckt p4_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p2_1
xr D G S B p2_1
.ends


* expanding   symbol:  n4_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n4_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n4_1.sch
.subckt n4_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n2_1
xl D G S B n2_1
.ends


* expanding   symbol:  p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_2.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  p2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p2_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p2_1.sch
.subckt p2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p1_1
xr D G S B p1_1
.ends


* expanding   symbol:  n2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n2_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n2_1.sch
.subckt n2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n1_1
xl D G S B n1_1
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_1.sym
* sch_path: /home/rodovalho/git/sky130amp/xschem/ampa/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
